module updown_counter (i_clk,
    i_rst,
    i_up_down,
    o_count);
 input i_clk;
 input i_rst;
 input i_up_down;
 output [3:0] o_count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net1;
 wire net2;

 INV_X1 _21_ (.A(net2),
    .ZN(_05_));
 AND2_X1 _22_ (.A1(_00_),
    .A2(_05_),
    .ZN(_01_));
 BUF_X2 _23_ (.A(net4),
    .Z(_06_));
 BUF_X4 _24_ (.A(i_up_down),
    .Z(_07_));
 XOR2_X1 _25_ (.A(_07_),
    .B(_00_),
    .Z(_08_));
 XNOR2_X1 _26_ (.A(_06_),
    .B(_08_),
    .ZN(_09_));
 NOR2_X1 _27_ (.A1(net2),
    .A2(_09_),
    .ZN(_02_));
 AND3_X1 _28_ (.A1(_06_),
    .A2(_07_),
    .A3(net3),
    .ZN(_10_));
 NOR3_X1 _29_ (.A1(_06_),
    .A2(_07_),
    .A3(net3),
    .ZN(_11_));
 OR3_X1 _30_ (.A1(net5),
    .A2(_10_),
    .A3(_11_),
    .ZN(_12_));
 OAI21_X1 _31_ (.A(net5),
    .B1(_10_),
    .B2(_11_),
    .ZN(_13_));
 AND3_X1 _32_ (.A1(_05_),
    .A2(_12_),
    .A3(_13_),
    .ZN(_03_));
 AND4_X1 _33_ (.A1(_06_),
    .A2(_07_),
    .A3(net5),
    .A4(net3),
    .ZN(_14_));
 NOR4_X1 _34_ (.A1(_06_),
    .A2(_07_),
    .A3(net5),
    .A4(net3),
    .ZN(_15_));
 OR3_X1 _35_ (.A1(net6),
    .A2(_14_),
    .A3(_15_),
    .ZN(_16_));
 OAI21_X1 _36_ (.A(net6),
    .B1(_14_),
    .B2(_15_),
    .ZN(_17_));
 AND3_X1 _37_ (.A1(_05_),
    .A2(_16_),
    .A3(_17_),
    .ZN(_04_));
 DFF_X1 \o_count[0]$_SDFF_PP0_  (.D(_01_),
    .CK(net1),
    .Q(net3),
    .QN(_00_));
 DFF_X1 \o_count[1]$_SDFF_PP0_  (.D(_02_),
    .CK(net1),
    .Q(net4),
    .QN(_20_));
 DFF_X1 \o_count[2]$_SDFF_PP0_  (.D(_03_),
    .CK(net1),
    .Q(net5),
    .QN(_19_));
 DFF_X1 \o_count[3]$_SDFF_PP0_  (.D(_04_),
    .CK(net1),
    .Q(net6),
    .QN(_18_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_47 ();
 BUF_X1 input1 (.A(i_clk),
    .Z(net1));
 BUF_X1 input2 (.A(i_rst),
    .Z(net2));
 BUF_X1 output3 (.A(net3),
    .Z(o_count[0]));
 BUF_X1 output4 (.A(net4),
    .Z(o_count[1]));
 BUF_X1 output5 (.A(net5),
    .Z(o_count[2]));
 BUF_X1 output6 (.A(net6),
    .Z(o_count[3]));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_73 ();
 FILLCELL_X32 FILLER_0_80 ();
 FILLCELL_X32 FILLER_0_112 ();
 FILLCELL_X32 FILLER_0_144 ();
 FILLCELL_X4 FILLER_0_176 ();
 FILLCELL_X2 FILLER_0_180 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X16 FILLER_1_161 ();
 FILLCELL_X4 FILLER_1_177 ();
 FILLCELL_X1 FILLER_1_181 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X16 FILLER_2_161 ();
 FILLCELL_X4 FILLER_2_177 ();
 FILLCELL_X1 FILLER_2_181 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X16 FILLER_3_161 ();
 FILLCELL_X4 FILLER_3_177 ();
 FILLCELL_X1 FILLER_3_181 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X16 FILLER_4_161 ();
 FILLCELL_X4 FILLER_4_177 ();
 FILLCELL_X1 FILLER_4_181 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X4 FILLER_5_73 ();
 FILLCELL_X32 FILLER_5_84 ();
 FILLCELL_X32 FILLER_5_116 ();
 FILLCELL_X32 FILLER_5_148 ();
 FILLCELL_X2 FILLER_5_180 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X16 FILLER_6_161 ();
 FILLCELL_X4 FILLER_6_177 ();
 FILLCELL_X1 FILLER_6_181 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_73 ();
 FILLCELL_X2 FILLER_7_77 ();
 FILLCELL_X1 FILLER_7_79 ();
 FILLCELL_X32 FILLER_7_84 ();
 FILLCELL_X32 FILLER_7_116 ();
 FILLCELL_X32 FILLER_7_148 ();
 FILLCELL_X2 FILLER_7_180 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_65 ();
 FILLCELL_X1 FILLER_8_73 ();
 FILLCELL_X16 FILLER_8_91 ();
 FILLCELL_X8 FILLER_8_107 ();
 FILLCELL_X2 FILLER_8_115 ();
 FILLCELL_X1 FILLER_8_117 ();
 FILLCELL_X4 FILLER_8_123 ();
 FILLCELL_X4 FILLER_8_132 ();
 FILLCELL_X4 FILLER_8_140 ();
 FILLCELL_X8 FILLER_8_149 ();
 FILLCELL_X4 FILLER_8_157 ();
 FILLCELL_X16 FILLER_8_164 ();
 FILLCELL_X2 FILLER_8_180 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_73 ();
 FILLCELL_X2 FILLER_9_77 ();
 FILLCELL_X1 FILLER_9_79 ();
 FILLCELL_X32 FILLER_9_86 ();
 FILLCELL_X4 FILLER_9_118 ();
 FILLCELL_X2 FILLER_9_122 ();
 FILLCELL_X1 FILLER_9_124 ();
 FILLCELL_X8 FILLER_9_129 ();
 FILLCELL_X4 FILLER_9_137 ();
 FILLCELL_X2 FILLER_9_141 ();
 FILLCELL_X1 FILLER_9_143 ();
 FILLCELL_X4 FILLER_9_161 ();
 FILLCELL_X2 FILLER_9_165 ();
 FILLCELL_X1 FILLER_9_167 ();
 FILLCELL_X8 FILLER_9_171 ();
 FILLCELL_X2 FILLER_9_179 ();
 FILLCELL_X1 FILLER_9_181 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_97 ();
 FILLCELL_X4 FILLER_10_113 ();
 FILLCELL_X2 FILLER_10_117 ();
 FILLCELL_X4 FILLER_10_124 ();
 FILLCELL_X32 FILLER_10_134 ();
 FILLCELL_X16 FILLER_10_166 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X16 FILLER_11_161 ();
 FILLCELL_X4 FILLER_11_177 ();
 FILLCELL_X1 FILLER_11_181 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X16 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_87 ();
 FILLCELL_X16 FILLER_12_119 ();
 FILLCELL_X4 FILLER_12_135 ();
 FILLCELL_X32 FILLER_12_144 ();
 FILLCELL_X4 FILLER_12_176 ();
 FILLCELL_X2 FILLER_12_180 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X8 FILLER_13_65 ();
 FILLCELL_X4 FILLER_13_73 ();
 FILLCELL_X32 FILLER_13_79 ();
 FILLCELL_X16 FILLER_13_111 ();
 FILLCELL_X8 FILLER_13_127 ();
 FILLCELL_X2 FILLER_13_135 ();
 FILLCELL_X1 FILLER_13_137 ();
 FILLCELL_X4 FILLER_13_142 ();
 FILLCELL_X16 FILLER_13_151 ();
 FILLCELL_X8 FILLER_13_167 ();
 FILLCELL_X4 FILLER_13_175 ();
 FILLCELL_X2 FILLER_13_179 ();
 FILLCELL_X1 FILLER_13_181 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_9 ();
 FILLCELL_X1 FILLER_14_11 ();
 FILLCELL_X32 FILLER_14_15 ();
 FILLCELL_X16 FILLER_14_47 ();
 FILLCELL_X8 FILLER_14_63 ();
 FILLCELL_X2 FILLER_14_71 ();
 FILLCELL_X4 FILLER_14_76 ();
 FILLCELL_X2 FILLER_14_80 ();
 FILLCELL_X1 FILLER_14_82 ();
 FILLCELL_X32 FILLER_14_87 ();
 FILLCELL_X32 FILLER_14_119 ();
 FILLCELL_X4 FILLER_14_151 ();
 FILLCELL_X1 FILLER_14_155 ();
 FILLCELL_X8 FILLER_14_173 ();
 FILLCELL_X1 FILLER_14_181 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X4 FILLER_15_65 ();
 FILLCELL_X1 FILLER_15_69 ();
 FILLCELL_X32 FILLER_15_87 ();
 FILLCELL_X32 FILLER_15_119 ();
 FILLCELL_X16 FILLER_15_151 ();
 FILLCELL_X8 FILLER_15_167 ();
 FILLCELL_X4 FILLER_15_178 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X16 FILLER_16_161 ();
 FILLCELL_X4 FILLER_16_177 ();
 FILLCELL_X1 FILLER_16_181 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X16 FILLER_17_161 ();
 FILLCELL_X4 FILLER_17_177 ();
 FILLCELL_X1 FILLER_17_181 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X16 FILLER_18_161 ();
 FILLCELL_X4 FILLER_18_177 ();
 FILLCELL_X1 FILLER_18_181 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X16 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_177 ();
 FILLCELL_X1 FILLER_19_181 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X16 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_177 ();
 FILLCELL_X1 FILLER_20_181 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X16 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_177 ();
 FILLCELL_X1 FILLER_21_181 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X4 FILLER_22_177 ();
 FILLCELL_X1 FILLER_22_181 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X8 FILLER_23_65 ();
 FILLCELL_X1 FILLER_23_73 ();
 FILLCELL_X32 FILLER_23_77 ();
 FILLCELL_X32 FILLER_23_109 ();
 FILLCELL_X32 FILLER_23_141 ();
 FILLCELL_X8 FILLER_23_173 ();
 FILLCELL_X1 FILLER_23_181 ();
endmodule
